module Shifter( dataA, dataB, dataOut );
input [31:0] dataA ;
input [4:0] dataB ;
output [31:0] dataOut ;

wire [31:0] layer1, layer2, layer3, layer4;
    // Layer 1: Shift by 1 bit
	mux mux0( .s(dataB[0]),.i0( 1'b0 ), .i1( dataA[0]), .o(layer1[0] ));
	mux mux1( .s(dataB[0]),.i0(dataA[0]), .i1( dataA[1]), .o(layer1[1] ));
	mux mux2( .s(dataB[0]),.i0(dataA[1]), .i1( dataA[2]), .o(layer1[2] ));
	mux mux3( .s(dataB[0]),.i0(dataA[2]), .i1( dataA[3]), .o(layer1[3] ));
	mux mux4( .s(dataB[0]),.i0(dataA[3]), .i1( dataA[4]), .o(layer1[4] ));
	mux mux5( .s(dataB[0]),.i0(dataA[4]), .i1( dataA[5]), .o(layer1[5] ));
	mux mux6( .s(dataB[0]),.i0(dataA[5]), .i1( dataA[6]), .o(layer1[6] ));
	mux mux7( .s( dataB[0]),.i0(dataA[6]), .i1( dataA[7]), .o(layer1[7] ));
	mux mux8( .s(dataB[0]),.i0(dataA[7]), .i1( dataA[8]), .o(layer1[8] ));
	mux mux9( .s(dataB[0]),.i0(dataA[8]), .i1( dataA[9]), .o(layer1[9] ));
	mux mux10( .s(dataB[0]),.i0(dataA[9]), .i1( dataA[10]), .o(layer1[10] ));
	mux mux11( .s(dataB[0]),.i0(dataA[10]), .i1( dataA[11]), .o(layer1[11] ));
	mux mux12( .s(dataB[0]),.i0(dataA[11]), .i1( dataA[12]), .o(layer1[12] ));
	mux mux13( .s(dataB[0]),.i0(dataA[12]), .i1( dataA[13]), .o(layer1[13] ));
	mux mux14( .s(dataB[0]),.i0(dataA[13]), .i1( dataA[14]), .o(layer1[14] ));
	mux mux15( .s(dataB[0]),.i0(dataA[14]), .i1( dataA[15]), .o(layer1[15] ));
	mux mux16( .s(dataB[0]),.i0(dataA[15]), .i1( dataA[16]), .o(layer1[16] ));
	mux mux17(.s( dataB[0]),.i0(dataA[16]), .i1( dataA[17]), .o(layer1[17] ));
	mux mux18( .s( dataB[0]),.i0(dataA[17]), .i1( dataA[18]), .o(layer1[18] ));
	mux mux19( .s(dataB[0]),.i0(dataA[18]), .i1( dataA[19]), .o(layer1[19] ));
	mux mux20( .s( dataB[0]),.i0(dataA[19]), .i1( dataA[20]), .o(layer1[20] ));
	mux mux21(  .s(dataB[0]),.i0(dataA[20]), .i1( dataA[21]), .o(layer1[21] ));
	mux mux22(  .s(dataB[0]),.i0(dataA[21]), .i1( dataA[22]), .o(layer1[22] ));
	mux mux23( .s( dataB[0]),.i0(dataA[22]), .i1( dataA[23]), .o(layer1[23] ));
	mux mux24( .s( dataB[0]),.i0(dataA[23]), .i1( dataA[24]), .o(layer1[24] ));
	mux mux25( .s( dataB[0]),.i0(dataA[24]), .i1( dataA[25]), .o(layer1[25] ));
	mux mux26( .s( dataB[0]),.i0(dataA[25]), .i1( dataA[26]), .o(layer1[26] ));
	mux mux27( .s( dataB[0]),.i0(dataA[26]), .i1( dataA[27]), .o(layer1[27] ));
	mux mux28( .s( dataB[0]),.i0(dataA[27]), .i1( dataA[28]), .o(layer1[28] ));
	mux mux29( .s( dataB[0]),.i0(dataA[28]), .i1( dataA[29]), .o(layer1[29] ));
	mux mux30( .s( dataB[0]),.i0(dataA[29]), .i1( dataA[30]), .o(layer1[30] ));
	mux mux31( .s( dataB[0]),.i0(dataA[30]), .i1( dataA[31]), .o(layer1[31] ));

    // Layer 3: Shift by 4 bits
	mux mux32( .s( dataB[1]),.i0( 1'b0), .i1(  layer1[0]), .o(layer2[0] ));
	mux mux33( .s( dataB[1]),.i0(1'b0), .i1( layer1[1]), .o(layer2[1] ));
	mux mux34( .s( dataB[1]),.i0(layer1[0]), .i1( layer1[2]), .o(layer2[2] ));
	mux mux35( .s( dataB[1]),.i0(layer1[1]), .i1( layer1[3]), .o(layer2[3] ));
	mux mux36( .s( dataB[1]),.i0(layer1[2]), .i1( layer1[4]), .o(layer2[4] ));
	mux mux37( .s( dataB[1]),.i0(layer1[3]), .i1( layer1[5]), .o(layer2[5] ));
	mux mux38( .s( dataB[1]),.i0(layer1[4]), .i1( layer1[6]), .o(layer2[6] ));
	mux mux39( .s( dataB[1]),.i0( layer1[5]), .i1( layer1[7]), .o(layer2[7] ));
	mux mux40( .s( dataB[1]),.i0(layer1[6]), .i1( layer1[8]), .o(layer2[8] ));
	mux mux41( .s( dataB[1]),.i0(layer1[7]), .i1( layer1[9]), .o(layer2[9] ));
	mux mux42( .s( dataB[1]),.i0( layer1[8]), .i1( layer1[10]), .o(layer2[10] ));
	mux mux43( .s( dataB[1]),.i0( layer1[9]), .i1( layer1[11]), .o(layer2[11] ));
	mux mux44( .s( dataB[1]),.i0( layer1[10]), .i1( layer1[12]), .o(layer2[12] ));
	mux mux45( .s( dataB[1]),.i0( layer1[11]), .i1( layer1[13]), .o(layer2[13] ));
	mux mux46( .s( dataB[1]),.i0( layer1[12]), .i1( layer1[14]), .o(layer2[14] ));
	mux mux47( .s( dataB[1]),.i0( layer1[13]), .i1( layer1[15]), .o(layer2[15] ));
	mux mux48( .s( dataB[1]),.i0( layer1[14]), .i1( layer1[16]), .o(layer2[16] ));
	mux mux49( .s( dataB[1]),.i0( layer1[15]), .i1( layer1[17]), .o(layer2[17] ));
	mux mux50( .s( dataB[1]),.i0( layer1[16]), .i1( layer1[18]), .o(layer2[18] ));
	mux mux51( .s( dataB[1]),.i0( layer1[17]), .i1( layer1[19]), .o(layer2[19] ));
	mux mux52( .s( dataB[1]),.i0( layer1[18]), .i1( layer1[20]), .o(layer2[20] ));
	mux mux53( .s( dataB[1]),.i0( layer1[19]), .i1( layer1[21]), .o(layer2[21] ));
	mux mux54( .s( dataB[1]),.i0( layer1[20]), .i1( layer1[22]), .o(layer2[22] ));
	mux mux55( .s( dataB[1]),.i0( layer1[21]), .i1( layer1[23]), .o(layer2[23] ));
	mux mux56( .s( dataB[1]),.i0( layer1[22]), .i1( layer1[24]), .o(layer2[24] ));
	mux mux57( .s( dataB[1]),.i0( layer1[23]), .i1( layer1[25]), .o(layer2[25] ));
	mux mux58( .s( dataB[1]),.i0( layer1[24]), .i1( layer1[26]), .o(layer2[26] ));
	mux mux59( .s(  dataB[1]),.i0( layer1[25]), .i1( layer1[27]), .o(layer2[27] ));
	mux mux60( .s( dataB[1]),.i0( layer1[26]), .i1( layer1[28]), .o(layer2[28] ));
	mux mux61( .s( dataB[1]),.i0( layer1[27]), .i1( layer1[29]), .o(layer2[29] ));
	mux mux62( .s( dataB[1]),.i0( layer1[28]), .i1( layer1[30]), .o(layer2[30] ));
	mux mux63( .s( dataB[1]),.i0( layer1[29]), .i1( layer1[31]), .o(layer2[31] ));

    // Layer 4: Shift by 8 bits
	mux mux64( .s( dataB[ 2]),.i0( 1'b0), .i1(layer2[0]), .o(layer3[ 0] ));
	mux mux65( .s(dataB[ 2]),.i0( 1'b0), .i1(layer2[1]), .o(layer3[ 1] ));
	mux mux66( .s(dataB[ 2]),.i0( 1'b0), .i1(layer2[2]), .o(layer3[ 2] ));
	mux mux67( .s(dataB[ 2]),.i0( 1'b0), .i1(layer2[3]), .o(layer3[ 3] ));
	mux mux68( .s(dataB[ 2]),.i0( layer2[0]), .i1(layer2[4]), .o(layer3[ 4] ));
	mux mux69(.s( dataB[ 2]),.i0( layer2[1]), .i1(layer2[5]), .o(layer3[ 5] ));
	mux mux70( .s(dataB[ 2]),.i0( layer2[2]), .i1(layer2[6]), .o(layer3[ 6] ));
	mux mux71(.s(dataB[ 2]),.i0( layer2[3]), .i1(layer2[7]), .o(layer3[ 7] ));
	mux mux72(.s(dataB[ 2]),.i0( layer2[4]), .i1(layer2[8]), .o(layer3[ 8] ));
	mux mux73(.s(dataB[ 2]),.i0( layer2[5]), .i1(layer2[9]), .o(layer3[ 9] ));
	mux mux74(.s(dataB[ 2]),.i0( layer2[6]), .i1(layer2[10]), .o(layer3[ 10] ));
	mux mux75(.s(dataB[ 2]),.i0( layer2[7]), .i1(layer2[11]), .o(layer3[ 11] ));
	mux mux76(.s(dataB[ 2]),.i0( layer2[8]), .i1(layer2[12]), .o(layer3[ 12] ));
	mux mux77(.s(dataB[ 2]),.i0( layer2[9]), .i1(layer2[13]), .o(layer3[ 13] ));
	mux mux78(.s(dataB[ 2]),.i0( layer2[10]), .i1(layer2[14]), .o(layer3[ 14] ));
	mux mux79(.s(dataB[ 2]),.i0( layer2[11]), .i1(layer2[15]), .o(layer3[ 15] ));
	mux mux80(.s(dataB[ 2]),.i0( layer2[12]), .i1(layer2[16]), .o(layer3[ 16] ));
	mux mux81(.s(dataB[ 2]),.i0( layer2[13]), .i1(layer2[17]), .o(layer3[ 17] ));
	mux mux82(.s(dataB[ 2]),.i0( layer2[14]), .i1(layer2[18]), .o(layer3[ 18] ));
	mux mux83(.s(dataB[ 2]),.i0( layer2[15]), .i1(layer2[19]), .o(layer3[ 19] ));
	mux mux84(.s(dataB[ 2]),.i0( layer2[16]), .i1(layer2[20]), .o(layer3[ 20] ));
	mux mux85(.s(dataB[ 2]),.i0( layer2[17]), .i1(layer2[21]), .o(layer3[ 21] ));
	mux mux86(.s(dataB[ 2]),.i0( layer2[18]), .i1(layer2[22]), .o(layer3[ 22] ));
	mux mux87(.s(dataB[ 2]),.i0( layer2[19]), .i1(layer2[23]), .o(layer3[ 23] ));
	mux mux88(.s(dataB[ 2]),.i0( layer2[20]), .i1(layer2[24]), .o(layer3[ 24] ));
	mux mux89(.s(dataB[ 2]),.i0( layer2[21]), .i1(layer2[25]), .o(layer3[ 25] ));
	mux mux90(.s(dataB[ 2]),.i0( layer2[22]), .i1(layer2[26]), .o(layer3[ 26] ));
	mux mux91(.s(dataB[ 2]),.i0( layer2[23]), .i1(layer2[27]), .o(layer3[ 27] ));
	mux mux92(.s(dataB[ 2]),.i0( layer2[24]), .i1(layer2[28]), .o(layer3[ 28] ));
	mux mux93(.s(dataB[ 2]),.i0( layer2[25]), .i1(layer2[29]), .o(layer3[ 29] ));
	mux mux94(.s(dataB[ 2]),.i0( layer2[26]), .i1(layer2[30]), .o(layer3[ 30] ));
	mux mux95(.s(dataB[ 2]),.i0( layer2[27]), .i1(layer2[31]), .o(layer3[ 31] ));

	mux mux96(.s(dataB[3]),.i0( 1'b0), .i1( layer3[0]), .o(layer4[0]  ));
	mux mux97(.s(dataB[3]),.i0(1'b0), .i1( layer3[1]), .o(layer4[1]  ));
	mux mux98(.s(dataB[3]),.i0(1'b0), .i1( layer3[2]), .o(layer4[2]  ));
	mux mux99(.s(dataB[3]),.i0(1'b0), .i1( layer3[3]), .o(layer4[3]  ));
	mux mux100(.s(dataB[3]),.i0(1'b0), .i1( layer3[4]), .o(layer4[4]  ));
	mux mux101(.s(dataB[3]),.i0(1'b0), .i1( layer3[5]), .o(layer4[5]  ));
	mux mux102(.s(dataB[3]),.i0(1'b0), .i1( layer3[6]), .o(layer4[6]  ));
	mux mux103(.s(dataB[3]),.i0(1'b0), .i1( layer3[7]), .o(layer4[7]  ));
	mux mux104(.s(dataB[3]),.i0(layer3[0]), .i1( layer3[8]), .o(layer4[8]  ));
	mux mux105(.s(dataB[3]),.i0(layer3[1]), .i1( layer3[9]), .o(layer4[9]  ));
	mux mux106(.s(dataB[3]),.i0(layer3[2]), .i1( layer3[10]), .o(layer4[10]  ));
	mux mux107(.s(dataB[3]),.i0(layer3[3]), .i1( layer3[11]), .o(layer4[11]  ));
	mux mux108(.s(dataB[3]),.i0(layer3[4]), .i1( layer3[12]), .o(layer4[12]  ));
	mux mux109(.s(dataB[3]),.i0(layer3[5]), .i1( layer3[13]), .o(layer4[13]  ));
	mux mux110(.s(dataB[3]),.i0(layer3[6]), .i1( layer3[14]), .o(layer4[14]  ));
	mux mux111(.s(dataB[3]),.i0(layer3[7]), .i1( layer3[15]), .o(layer4[15]  ));
	mux mux112(.s(dataB[3]),.i0(layer3[8]), .i1( layer3[16]), .o(layer4[16]  ));
	mux mux113(.s(dataB[3]),.i0(layer3[9]), .i1( layer3[17]), .o(layer4[17]  ));
	mux mux114(.s(dataB[3]),.i0(layer3[10]), .i1( layer3[18]), .o(layer4[18]  ));
	mux mux115(.s(dataB[3]),.i0(layer3[11]), .i1( layer3[19]), .o(layer4[19]  ));
	mux mux116(.s(dataB[3]),.i0(layer3[12]), .i1( layer3[20]), .o(layer4[20]  ));
	mux mux117(.s(dataB[3]),.i0(layer3[13]), .i1( layer3[21]), .o(layer4[21]  ));
	mux mux118(.s(dataB[3]),.i0(layer3[14]), .i1( layer3[22]), .o(layer4[22]  ));
	mux mux119(.s(dataB[3]),.i0(layer3[15]), .i1( layer3[23]), .o(layer4[23]  ));
	mux mux120(.s(dataB[3]),.i0(layer3[16]), .i1( layer3[24]), .o(layer4[24]  ));
	mux mux121(.s(dataB[3]),.i0(layer3[17]), .i1( layer3[25]), .o(layer4[25]  ));
	mux mux122(.s(dataB[3]),.i0(layer3[18]), .i1( layer3[26]), .o(layer4[26]  ));
	mux mux123(.s(dataB[3]),.i0(layer3[19]), .i1( layer3[27]), .o(layer4[27]  ));
	mux mux124(.s(dataB[3]),.i0(layer3[20]), .i1( layer3[28]), .o(layer4[28]  ));
	mux mux125(.s(dataB[3]),.i0(layer3[21]), .i1( layer3[29]), .o(layer4[29]  ));
	mux mux126(.s(dataB[3]),.i0(layer3[22]), .i1( layer3[30]), .o(layer4[30]  ));
	mux mux127(.s(dataB[3]),.i0(layer3[23]), .i1( layer3[31]), .o(layer4[31]  ));
	
    // Layer 5: Shift by 16 bits
	mux mux128(.s(dataB[4]),.i0(1'b0), .i1( layer4[0]), .o(dataOut[0]  ));
	mux mux129(.s(dataB[4]),.i0(1'b0), .i1( layer4[1]), .o(dataOut[1]  ));
	mux mux130(.s(dataB[4]),.i0(1'b0), .i1( layer4[2]), .o(dataOut[2]  ));
	mux mux131(.s(dataB[4]),.i0(1'b0), .i1( layer4[3]), .o(dataOut[3]  ));
	mux mux132(.s(dataB[4]),.i0(1'b0), .i1( layer4[4]), .o(dataOut[4]  ));
	mux mux133(.s(dataB[4]),.i0(1'b0), .i1( layer4[5]), .o(dataOut[5]  ));
	mux mux134(.s(dataB[4]),.i0(1'b0), .i1( layer4[6]), .o(dataOut[6]  ));
	mux mux135(.s(dataB[4]),.i0(1'b0), .i1( layer4[7]), .o(dataOut[7]  ));
	mux mux136(.s(dataB[4]),.i0(1'b0), .i1( layer4[8]), .o(dataOut[8]  ));
	mux mux137(.s(dataB[4]),.i0(1'b0), .i1( layer4[9]), .o(dataOut[9]  ));
	mux mux138(.s(dataB[4]),.i0(1'b0), .i1( layer4[10]), .o(dataOut[10]  ));
	mux mux139(.s(dataB[4]),.i0(1'b0), .i1( layer4[11]), .o(dataOut[11]  ));
	mux mux140(.s(dataB[4]),.i0(1'b0), .i1( layer4[12]), .o(dataOut[12]  ));
	mux mux141(.s(dataB[4]),.i0(1'b0), .i1( layer4[13]), .o(dataOut[13]  ));
	mux mux142(.s(dataB[4]),.i0(1'b0), .i1( layer4[14]), .o(dataOut[14]  ));
	mux mux143(.s(dataB[4]),.i0(1'b0), .i1( layer4[15]), .o(dataOut[15]  ));
	mux mux144(.s(dataB[4]),.i0(layer4[0]), .i1( layer4[16]), .o(dataOut[16]  ));
	mux mux145(.s(dataB[4]),.i0(layer4[1]), .i1( layer4[17]), .o(dataOut[17]  ));
	mux mux146(.s(dataB[4]),.i0(layer4[2]), .i1( layer4[18]), .o(dataOut[18]  ));
	mux mux147(.s(dataB[4]),.i0(layer4[3]), .i1( layer4[19]), .o(dataOut[19]  ));
	mux mux148(.s(dataB[4]),.i0(layer4[4]), .i1( layer4[20]), .o(dataOut[20]  ));
	mux mux149(.s(dataB[4]),.i0(layer4[5]), .i1( layer4[21]), .o(dataOut[21]  ));
	mux mux150(.s(dataB[4]),.i0(layer4[6]), .i1( layer4[22]), .o(dataOut[22]  ));	
	mux mux151(.s(dataB[4]),.i0(layer4[7]), .i1( layer4[23]), .o(dataOut[23]  ));
	mux mux152(.s(dataB[4]),.i0(layer4[8]), .i1( layer4[24]), .o(dataOut[24]  ));
	mux mux153(.s(dataB[4]),.i0(layer4[9]), .i1( layer4[25]), .o(dataOut[25]  ));
	mux mux154(.s(dataB[4]),.i0(layer4[10]), .i1( layer4[26]), .o(dataOut[26]  ));
	mux mux155(.s(dataB[4]),.i0(layer4[11]), .i1( layer4[27]), .o(dataOut[27]  ));
	mux mux156(.s(dataB[4]),.i0(layer4[12]), .i1( layer4[28]), .o( dataOut[28]  ));
	mux mux157(.s(dataB[4]),.i0(layer4[13]), .i1( layer4[29]), .o( dataOut[29]  ));
	mux mux158(.s(dataB[4]),.i0(layer4[14]), .i1( layer4[30]), .o( dataOut[30]  ));	
	mux mux159(.s(dataB[4]),.i0(layer4[15]), .i1( layer4[31]), .o(dataOut[31]  ));
	


	
endmodule